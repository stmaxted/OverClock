
module InternalOsciallator (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
